-----------�ӵ�Ƭ�����յ�������DDSģ���������Ƶ���ֺ���λ������
-----------ռ�ձȿ�����
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
entity fifo_control is
port(
    f:in std_logic;--Ƶ��
    -- p:in std_logic;--��λ
    --h:in std_logic;--ռ�ձ�
    mcu_datain:in std_logic_vector(7 downto 0);--��Ƭ����������
    data_outf:out std_logic_vector(7 downto 0);---FIFO�������--Ƶ�ʿ���
    data_outh:out std_logic_vector(7 downto 0);--ռ�ձȿ�����
    w_req:in std_logic;--д����
    clk:in std_logic--ͬ��ʱ��
);
end fifo_control;
architecture behave of fifo_control is
---------------FIFO����------------------
component fifo_mcu
port(
     data:in std_logic_vector(7 downto 0);
     wrreq:in std_logic;
     rdreq:in std_logic;
     clock:in std_logic;
     q:out std_logic_vector(7 downto 0);
     full:out std_logic;
     empty:out std_logic
);
end component;
signal full_flag:std_logic;--����־
signal empty_flag:std_logic;--�ձ�־
signal clk_div:std_logic;--��Ƶ��ΪFIFO�Ĳ���ʱ��
signal r_req:std_logic;--������
signal data_temp:std_logic_vector(7 downto 0);
signal data_temp1:std_logic_vector(7 downto 0);
signal flag1,flag2:std_logic;
begin 
  u1: fifo_mcu port map(data=>mcu_datain,wrreq=>w_req,rdreq=>r_req,clock=>clk_div,q=>data_temp,full=>full_flag,empty=>empty_flag);
---------------��Ƶ(1MHz)------------------ 
 process(clk)
   variable counter:integer range 0 to 24;
    begin 
      if(clk'event and clk='1')then 
         if(counter=24)then 
             counter:=0;
         else 
             counter:=counter+1;
             clk_div<=not clk_div;
         end if;
      end if;
 end process;
 ------------------------------------
 data_temp1<=data_temp;
 ----------fifo������----------------
 process(f,empty_flag)
 begin
   if(f='1')then--Ƶ�ʱ�־
      if(empty_flag='0')then --δ�ձ�־
           r_req<='1';--������
           
         if(data_temp1="10000001")then--���ݷ���
               flag1<='1';
               flag2<='0;
         elsif(data_temp="01000010")then--���ݷ���
               flag2<='1';
               flag1<='0';
         else null;
         end if;    
      else
          null;
      end if;
   end if;
 end process;
 process(flag1,flag2,clk)
    begin 
      if(clk'event and clk='1')then 
          if(flag1='1')then 
              data_outf<=data_temp1;--Ƶ��
          end if;
          if(flag2='1')then
              data_outh<=data_temp1;--ռ�ձ�
          end if;
      end if;
 end process;  
end behave;





