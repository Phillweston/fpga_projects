/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� DDS_top.v
** �������ڣ�
** �����������������
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module DDS_top(clk,                                 //�ڲ�ʱ��
               reset,                               //��λ�ź� key5
               sclk,                                //TLC5615 sclkʱ�ӽ�
               din,                                 //TLC5615 din���ݽ�
               cs,                                  //TLC5615 csƬѡ
               set_waveform_key_in,                 //�������ð��� key1
               set_f_key_in,                        //Ƶ�����ð��� key2
               set_a_key_in,                        //��ֵ���ð��� key3
               set_p_key_in,                        //��λ���ð��� key4
               sin_data                             //����Ĳ������ݣ����ڲ���
              );
input      clk;
input      reset;
input      set_waveform_key_in;
input      set_f_key_in,set_a_key_in,set_p_key_in;
output     din;
output     cs;
output     sclk;
output     [9:0]sin_data;

wire clk;
wire reset;
wire set_waveform_key_in;
wire set_f_key_in,set_a_key_in,set_p_key_in;

wire [1:0] set_waveform_line;
wire [20:0] f_control_line;
wire [3:0]  a_control_line;
wire [8:0]  p_control_line;

wire       set_waveform_key;
wire       set_f_key;
wire       set_a_key;
wire       set_p_key;
//ģ������
    //DDsģ��
  DDS     u4(
             .clk(clk),
             .dds_data_out(sin_data),
             .set_waveform(set_waveform_line),
             .set_f(f_control_line),
             .set_a(a_control_line),
             .set_p(p_control_line)
             );
    //DAC����ģ��
  TLC5615 U5(.clk(clk),.sclk(sclk),.din(din),.cs(cs),.din_in(sin_data));
    //��������ģ��
  key     u6(.clk(clk),.key(set_waveform_key_in),.key_out(set_waveform_key));
  key     u7(.clk(clk),.key(set_f_key_in),.key_out(set_f_key));
  key     u8(.clk(clk),.key(set_a_key_in),.key_out(set_a_key));
  key     u9(.clk(clk),.key(set_p_key_in),.key_out(set_p_key));
    //��������ģ��
  key_coding u10(
                .reset(reset),
                .set_waveform_key(set_waveform_key),
                .set_f_key(set_f_key),
                .set_a_key(set_a_key),
                .set_p_key(set_p_key),
                .set_waveform(set_waveform_line),
                .f_control(f_control_line),
                .a_control(a_control_line),
                .p_control(p_control_line));

endmodule


