-- ******************************************************************************
-- ����ģ��
-- *******************************************************************************
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
entity control is
port(
    clk:in std_logic;                               --50Mʱ������
    reset_n:in std_logic;                           --��λ�ź�����
    start_signal:in std_logic;                      --��ʼ����
    mileage_signal:in std_logic;                    --��̰�����ÿ��һ���������1����
    wait_signal:in std_logic;                       --�ȴ�����
    
    mileage_counter_ge_out:out std_logic_vector(3 downto 0);
    mileage_counter_shi_out:out std_logic_vector(3 downto 0);
    
    
    minute_out:out integer range 60 downto 0;       --����ȴ���������
    mileage_out:out integer range 99 downto 0;      --�����ʻ������
    cost_out:out integer range 99 downto 0         --�������
);
end control;
architecture control_behave of control is 
type state is(
            prepare_state,--׼��״̬
            start_state,--��ʼ״̬
            wait_state,--�ȴ�״̬
            arrive_state--�������״̬
            );
signal  current_state:state;--һ��ʼ����׼��״̬
signal  start_flag:std_logic;--������ʼ�źű�־
signal  wait_flag:std_logic_vector(1 downto 0);--�����ȴ��źű�־
signal  mileage_counter:integer range 99 downto 0;--��¼��ʻ������
signal  mileage_counter_ge:std_logic_vector(3 downto 0);
signal  mileage_counter_shi:std_logic_vector(3 downto 0);
signal  cost_counter:integer range 99 downto 0;
signal  cost_counter_temp1:integer range 99 downto 0;
signal  cost_counter_temp2:integer range 99 downto 0;
signal  temp1:integer range 99 downto 0;
signal  temp2:integer range 99 downto 0;
signal  temp3:integer range 99 downto 0;
signal  minute_counter:integer range 60 downto 0;
signal  count:integer range 250000 downto 0;--��Ƶ������
signal  second_count:integer range 6000 downto 0;--�������
signal  clk_div:std_logic; --��Ƶʱ��
begin
    --������á���̡����ӵ�����
    minute_out <= minute_counter;
    mileage_out <= mileage_counter;
    mileage_counter_ge_out <= mileage_counter_ge;
    mileage_counter_shi_out <= mileage_counter_shi;
    cost_out <= cost_counter;
    
    -- //****************************************************************************************************
    -- //  ģ������:��ʼ�������ģ�飬�����¿�ʼ�������൱����������
    -- //  ��������:start_flagΪ��1��ʱ����ʾ��ʼ
    -- //****************************************************************************************************
    process(start_signal,reset_n)
    begin
        if(reset_n = '0')then
            start_flag <= '0';
        elsif(start_signal'event and start_signal = '0')then--�½��ش���
            start_flag <= '1';
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:��̰���������ʻ��������ÿ��һ�Σ�����������1����
    -- //  ��������:
    -- //****************************************************************************************************
    process(mileage_signal,reset_n)
    begin
        if(reset_n = '0')then
            mileage_counter <= 0;
        elsif(mileage_signal'event and mileage_signal = '0')then--�½��ش���
            if(start_flag = '1')then
                if(mileage_counter = 99)then
                    mileage_counter <= 0;
                else
                    mileage_counter <= mileage_counter + 1;
                end if;
            end if;
        end if;
    end process;
    process(mileage_signal,reset_n)
    begin
        if(reset_n = '0')then
            mileage_counter_ge <= "0000";
            mileage_counter_shi <= "0000";
        elsif(mileage_signal'event and mileage_signal = '0')then
            if(start_flag = '1')then
                if(mileage_signal = '0')then--����������
                    if(mileage_counter_ge = "1001")then
                        if(mileage_counter_shi = "1001")then
                            mileage_counter_shi <= "0000";
                        else
                            mileage_counter_ge <= "0000";
                            mileage_counter_shi <= mileage_counter_shi + '1';
                        end if;
                    else
                        mileage_counter_ge <= mileage_counter_ge + '1';
                    end if;
                end if;
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:�ȴ���������һ�ΰ��µȴ�������ͣ���ȴ�������ȴ���ʱ״̬���ٰ�һ�Σ��˳��ȴ���ʱ״̬
    -- //  ��������:wait_flagΪ��1��ʱ����ʾ��ʼ
    -- //****************************************************************************************************
    process(wait_signal,reset_n)
    begin
        if(reset_n = '0')then
            wait_flag <= "00";
        elsif(wait_signal'event and wait_signal = '0')then--�½��ش���
            if(wait_flag = "00")then
                wait_flag <= "01";--��01���ȴ���־
            else
                wait_flag <= not wait_flag;--����ȡ��
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:��Ƶģ��
    -- //  ��������:��50Mʱ�ӷ���100Hz
    -- //****************************************************************************************************
    process(clk,reset_n)--100HZ
      begin 
        if(reset_n = '0')then
            count <= 0;
            clk_div <= '0';
        elsif(clk'event and clk = '1')then--�����ش���
            if(count = 249999)then--
                count <= 0;
                clk_div <= not clk_div;
            else
                count <= count + 1;
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:���ʱģ��
    -- //  ��������:��100Hz�������ʱ
    -- //****************************************************************************************************
    process(clk,reset_n)--100HZ
      begin 
        if(reset_n = '0')then
            second_count <= 0;
            minute_counter <= 0;
        elsif(clk'event and clk = '1')then--�����ش���
            if(start_flag = '1')then
                if(wait_flag = "01")then--����ȴ�״̬�Ž��м�ʱ
                    if(second_count = 6000)then--
                        second_count <= 0;
                        if(minute_counter = 60)then
                            minute_counter <= 0;
                        else
                            minute_counter <= minute_counter + 1;
                        end if;
                    else
                        second_count <= second_count + 1;
                    end if;
                 end if;
             end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:�������
    -- //  ��������:
    -- //****************************************************************************************************
    temp1 <= mileage_counter - 3;
    temp2 <= temp1 * 2;
    cost_counter_temp1 <= 6 + temp2 + minute_counter;
    
    temp3 <= mileage_counter * 2;
    cost_counter_temp2 <= temp3 + minute_counter;

    process(clk_div,reset_n)
    begin
        if(reset_n = '0')then
            cost_counter <= 0;
        elsif(clk_div'event and clk_div = '1')then--
            if(start_flag = '1')then
                if(mileage_counter <= 3)then--������С�ڻ��ߵ���3����
                    cost_counter <= 6;
                elsif(mileage_counter > 3 and mileage_counter <= 19)then--����������3���С�ڻ��ߵ���19����
                    cost_counter <= cost_counter_temp1;
                elsif(mileage_counter > 19)then--����������3���С�ڻ��ߵ���19����
                    cost_counter <= cost_counter_temp2;
                else--����������19����
                    NULL;
                end if;
            end if;
        end if;
    end process;

end control_behave;












