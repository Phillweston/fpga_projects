----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    
-- Design Name: 
-- Module Name:    enemy - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--������ʾ����ʾ���ķɻ���״���ã�������ַ���0��ɵľ��Ƿɻ���ģ��
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity enemy is
    port(
        y,x: in std_logic_vector(5 downto 0);----location of point��y����ĳһ�У�x����ĳһ�У����Ƕ�ά����
        data: out std_logic---yan se xin xi�ɻ�����ɫ�ź�
    );
end enemy;

architecture Behavioral of enemy is
    type rom_type is array(0 to 31) of std_logic_vector(31 downto 0);
    constant FONT: rom_type :=
    ("11111111111111111111111111111111",
     "11111111100001100110000111111111",
     "11111111111000111100011111111111",
     "11111111111110000001111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111110011001111111111111",
     "11111111111110011001111111111111",
     "11000000111110000001111100000011",
     "11000000001110000001110000000011",
     "11001101000000111100000010110011",
     "11111101110000100100001110111111",
     "11111101111100000000111110111111",
     "11111101111111100001111110111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111110000001111111111111",
     "11111111111111000011111111111111",
     "11111111111111100111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111");

signal d:std_logic_vector(31 downto 0);
begin 

d<=FONT(conv_integer(y));
data<=not d(conv_integer(x));

end Behavioral;

