----------------------------------------------------------------------
----------------------------------------------------------------------
-- (�������ݵĹ���)��ʼ����׼�������ʹӻ���ַ������Ӧ��
--                  �����ֽڵ�ַ������Ӧ�𣬷������ݣ�����Ӧ��
--                  ����ֹͣ�ź�
----------------------------------------------------------------------
-- (�������ݵĹ���)��ʼ����׼�������ʹӻ���ַ������Ӧ��
--                  �����ֽڵ�ַ������Ӧ��
----------------------------------------------------------------------
-- ��ʼ��1�����ʹӻ���ַ������Ӧ�𣬶�ȡ���ݣ�����ֹͣ�źţ�����״̬
----------------------------------------------------------------------
-- ��д���������ú󣬽��ж�����
----------------------------------------------------------------------
-- �������ã�scl��24��sda��26
-- 4�������ֱ�Ϊ��74��67��70��72
-- 4��LED�ֱ�Ϊ��141��142��143��144
----------------------------------------------------------------------
-- ����˵����ͨ���������������ʽ���沦�뿪�صĹ���
----------------------------------------------------------------------
-- key1Ϊȷ�ϰ�����ÿ���Ȱ���key2~key5�İ�����Ȼ����key1�������ͽ�������
--      ��Ϣͨ��iic���͵�iicоƬ��AT24c04���ϣ�Ȼ�������ʾ��led��
----------------------------------------------------------------------
-- key2Ϊ��ͨ����������Ϊ0������Ϊ1����Ӧled4�����²��ſ���ͬʱ����key1��ſ�����
--      �����ݡ�0111��ͨ��iic���͵�iicоƬ����ͨ��iic������ʾ��led�ϣ���ʱ��led4��������LED������
----------------------------------------------------------------------
-- key3Ϊ��ͨ����������Ϊ0������Ϊ1����Ӧled3�����²��ſ���ͬʱ����key1��ſ�����
--      �����ݡ�1011��ͨ��iic���͵�iicоƬ����ͨ��iic������ʾ��led�ϣ���ʱ��led3��������LED������
----------------------------------------------------------------------
-- key4Ϊ��ͨ����������Ϊ0������Ϊ1����Ӧled2�����²��ſ���ͬʱ����key1��ſ�����
--      �����ݡ�1101��ͨ��iic���͵�iicоƬ����ͨ��iic������ʾ��led�ϣ���ʱ��led2��������LED������
----------------------------------------------------------------------
-- key5Ϊ��ͨ����������Ϊ0������Ϊ1����Ӧled1�����²��ſ���ͬʱ����key1��ſ�����
--      �����ݡ�1110��ͨ��iic���͵�iicоƬ����ͨ��iic������ʾ��led�ϣ���ʱ��led1��������LED������
----------------------------------------------------------------------
----------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
entity iic is
port(
    clk:in      std_logic;--�����50Mʱ���ź�
    reset_n:in  std_logic;--
    sda:inout   std_logic;--IIC�������ź�
    scl:inout   std_logic;--IIC��ʱ���ź�
    key:in      std_logic_vector(3 downto 0);       --��������
    led:out     std_logic_vector(7 downto 0);       --LED��ʾ�ź�
    seg_duan:out std_logic_vector(7 downto 0);      --����ܶ��ź����
    seg_wei:out std_logic_vector(7 downto 0)        --�����λ�ź����
);
end iic ;
architecture behave of iic  is
signal clk_div: std_logic;--��Ƶ���ʱ��

type state is(
            prepare,--׼��״̬
            start,--��ʼ״̬
            send_slave_address,--���ʹӻ���ַ״̬
            ask1,--Ӧ��״̬1
            send_bit_address,--���ʹ洢��ַ״̬
            ask2,--Ӧ��״̬2
            send_data,--��������
            nack,--û��Ӧ��״̬
            start1,--��ʼ״̬
            send_read,--����Ҫ���ж�����״̬
            ask3,--Ӧ��״̬3
            read_data,--��ȡ����
            stop,--����
            idle--����״̬
            );
signal current_state:state := prepare;--һ��ʼ����׼��״̬
signal slave_address:   std_logic_vector(8 downto 1):="10100000";--�ӻ���ַ
signal bit_address:     std_logic_vector(8 downto 1):="00000001";--�ֽڵ�ַ
signal data:            std_logic_vector(8 downto 1):="11110000";---�����͵�����
signal data_temp:       std_logic_vector(8 downto 1);--�������ݼĴ���
signal flag_rw:         std_logic:='0';             --��дת����־
signal clk_1hz:         std_logic;
signal count:           std_logic_vector(24 downto 0);
signal clk_scan:        std_logic;
signal seg_select:      std_logic_vector(1 downto 0);
signal scan_count:      std_logic_vector(13 downto 0);
signal data_temp_shi:   std_logic_vector(3 downto 0);
signal data_temp_ge:    std_logic_vector(3 downto 0);
begin
    ----------------------------------------------------------------------
    -- ��Ƶ��������50Mʱ�ӷ�Ƶ��1KHz
    ----------------------------------------------------------------------
    process(clk)
    variable counter:   integer range 0 to 25000;
    begin 
        if(clk'event and clk = '1')then  
            if(counter = 24999)then 
                counter := 0;
                clk_div <= not clk_div;
            else 
                counter := counter + 1;
            end if;
        end if;
    end process;
    ----------------------------------------------------------------------
    -- ��������״̬�ɼ���������������״̬Ϊ��1������Ӧ��led����û�а���״̬Ϊ��0������Ӧ��led��
    ----------------------------------------------------------------------
    ----------------------------------------------------------------------
    -- iicͨ��д�������ģ��
    ----------------------------------------------------------------------
    process(clk_div,reset_n)
    variable counter:       integer range 0 to 20;
    variable num_counter:   integer range 0 to 8:=8;--�������ݼ����Ĵ���
    variable temp:          std_logic_vector(6 downto 0);
    begin 
        if(reset_n = '0')then
            led <= "11111111";--led��
            --��������״̬�ɼ���������������״̬Ϊ��1������Ӧ��led����û�а���״̬Ϊ��0������Ӧ��led��
            data(4 downto 1) <= key(3 downto 0);
            
            slave_address(8 downto 1)<="10100000";--�ӻ���ַ
            bit_address(8 downto 1)<="00000001";--�ֽڵ�ַ
            current_state <= prepare;--׼��״̬
            num_counter:=8;
            counter:=0;
            temp:="0000000";
            flag_rw<='0';
        elsif(clk_div'event and clk_div = '1')then 
    --------------------------------------------
    --------------------����д��״̬-----------
    --------------------------------------------
            if(flag_rw = '0')then
                case current_state is
                    when prepare=>temp:=temp+1;---����׼��״̬
                        if(temp="0000010")then 
                            temp:="0000000";
                            current_state<=start;
                        else
                            current_state<=prepare;
                        end if;
                    when start=>---������ʼ�ź�
                        counter:=counter+1;
                        case counter is
                            when 1=>sda<='1';
                            when 2=>scl<='1';
                            when 3=>sda<='0';
                            when 4=>scl<='0';
                            when 5=>counter:=0;
                            current_state<=send_slave_address;
                            when others=>null;
                        end case;
                    when send_slave_address=>--���ʹӻ���ַ
                        counter:=counter+1;
                        -- led<="01111111";
                        case counter is
                            when 1=>sda<=slave_address(num_counter);---�ȷ��͸�λ����
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then--�ж�8λ�����Ƿ�����
                                    current_state<=ask1;
                                    num_counter:=8;
                                else 
                                    current_state<=send_slave_address;
                                end if;
                            when others=>null;
                        end case;
                    when ask1=>--Ӧ��1
                        counter:=counter+1;
                        -- led<="10111111";
                        case counter is
                            when 1=>sda<='0';
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>counter:=0;
                                current_state<=send_bit_address;
                            when others=>null;
                        end case;
                    when send_bit_address=>--�����ֽڵ�ַ
                        counter:=counter+1;
                        -- led<="11011111";
                        case counter is
                            when 1=>sda<=bit_address(num_counter);
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>
                                num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then 
                                    current_state<=ask2;
                                    num_counter:=8;
                                else 
                                    current_state<=send_bit_address;
                                end if;
                            when others=>null;
                        end case;
                    when ask2=>counter:=counter+1;---Ӧ��2
                        -- led<="11101111";
                        case counter is
                            when 1=>sda<='0';
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>counter:=0;
                            current_state<=send_data;
                            when others=>null;
                        end case;
                    when send_data=>counter:=counter+1;--��������
                        -- led<="11110111";
                        case counter is
                            when 1=>sda<=data(num_counter);
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>
                                num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then 
                                    current_state<=ask3;
                                    num_counter:=8;
                                else 
                                    current_state<=send_data;
                                end if;
                            when others=>null;
                        end case;
                    when ask3=>--Ӧ��3
                        counter:=counter+1;
                        -- led<="11111011";
                        case counter is
                            when 1=>sda<='0';
                            when 2=>scl<='1';
                            when 3=>scl<='0';
                            when 4=>counter:=0;
                                current_state<=stop;
                            when others=>null;
                        end case;
                    when stop=>--ֹͣ�ź�
                        counter:=counter+1;
                        -- led<="11111101";
                        case counter is
                            when 1=>sda<='0';
                            when 3=>scl<='1';
                            when 10=>sda<='1';
                            when 15=>counter:=0;
                            current_state<=idle;
                            when others=>null;
                        end case;
                    when idle=>sda<='1';---����
                        scl<='1';
                        current_state<=prepare;
                        -- led<="11111110";
                        flag_rw<='1';--״̬ת������ȡ����
                        ---��ʼ��
                        num_counter:=8;
                        counter:=0;
                        temp:="0000000";
                        when others=>null;
                end case;
            end if;
    ------------------------------------------------------
    ----------------�����ȡ״̬-------------------------
    ------------------------------------------------------
            if(flag_rw = '1')then
                case current_state is
                    when prepare=>temp:=temp+1;
                        if(temp="0000010")then 
                            temp:="0000000";
                            current_state<=start;
                        else
                            current_state<=prepare;
                        end if;
                    when start=>
                        counter:=counter+1;
                        case counter is
                            when 1=>sda<='1';
                            when 3=>scl<='1';
                            when 5=>sda<='0';
                            when 7=>scl<='0';
                            when 9=>counter:=0;
                                current_state<=send_slave_address;
                            when others=>null;
                        end case;
                    when send_slave_address=>
                        counter:=counter+1;
                        -- led<="01111111";
                        case counter is
                            when 1=>sda<=slave_address(num_counter);---�ȷ��͸�λ����
                            when 3=>scl<='1';
                            when 6=>scl<='0';
                            when 8=>num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then--�ж�8λ�����Ƿ�����
                                    current_state<=ask1;
                                    num_counter:=8;
                                else 
                                    current_state<=send_slave_address;
                                end if;
                            when others=>null;
                        end case;    
                    when ask1=>
                        counter:=counter+1;
                        -- led<="10111111";
                        case counter is
                            when 3=>sda<='0';
                            when 6=>scl<='1';
                            when 8=>scl<='0';
                            when 10=>counter:=0;
                                current_state<=send_bit_address;
                            when others=>null;
                        end case;
                    when send_bit_address=>
                        counter:=counter+1;
                        -- led<="11011111";
                        case counter is
                            when 1=>sda<=bit_address(num_counter);
                            when 3=>scl<='1';
                            when 6=>scl<='0';
                            when 9=>
                                num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then 
                                    current_state<=ask2;
                                    num_counter:=8;
                                else 
                                    current_state<=send_bit_address;
                                end if;
                            when others=>null;
                        end case;
                    when ask2=>counter:=counter+1;
                        -- led<="11101111";
                        case counter is
                            when 3=>sda<='0';
                            when 6=>scl<='1';
                            when 8=>scl<='0';
                            when 10=>counter:=0;
                                current_state<=start1;
                            when others=>null;
                        end case;
                    when start1=>--���³�ʼ��
                        counter:=counter+1;
                        -- led<="11110111";
                        case counter is
                            when 1=>sda<='1';
                            when 3=>scl<='1';
                            when 6=>sda<='0';
                            when 8=>scl<='0';
                            when 10=>counter:=0;
                                current_state<=send_read;
                                slave_address<="10100001";
                            when others=>null;
                        end case;       
                    when send_read=>--���ʹӻ���ַ
                        counter:=counter+1;
                        -- led<="11111011";
                        case counter is
                            when 1=>sda<=slave_address(num_counter);
                            when 4=>scl<='1';
                            when 6=>scl<='0';
                            when 9=>num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then 
                                    num_counter:=8;
                                    current_state<=ask3;
                                else 
                                    current_state<=send_read;
                                end if;
                            when others=>null;
                        end case;
                    when ask3=>counter:=counter+1;--Ӧ��
                        -- led<="11111101";
                        case counter is
                            when 3=>sda<='0';
                            when 6=>scl<='1';
                            when 8=>scl<='0';
                            when 10=>current_state<=read_data;
                                counter:=0;
                            when others=>null;
                            end case;
                    when read_data=>--��ȡ����
                        counter:=counter+1;
                        -- led<="11111110";
                        case counter is
                            when 1=>sda<='Z';
                            when 4=>scl<='1';
                            when 8=>data_temp(num_counter)<=sda;
                            when 10=>scl<='0';
                            when 12=>num_counter:=num_counter-1;
                                counter:=0;
                                if(num_counter=0)then 
                                    num_counter:=8;
                                    current_state<=stop;
                                else 
                                    current_state<=read_data;
                                end if;
                            when others=>null;
                        end case;
                        --ֹͣ�ź�(�ڶ�ȡһ������֮���������û��Ӧ���򣬴ӻ���AT24c04�����ڵȴ�״̬��
                        --����������һ��ֹͣ�źţ��ӻ����ڱ��õ�Դ״̬��)�����������Ӧ����ӻ�������������
                    when stop=>
                        counter:=counter+1;
                        case counter is
                            when 1=>sda<='0';
                            when 3=>scl<='1';
                            when 6=>sda<='1';
                            when 8=>counter:=0;
                                current_state<=idle;
                            when others=>null;
                        end case;
                    when idle=>sda<='1';--����
                        scl<='1';
                        led<=data_temp;
                        current_state <= idle;--���½���д����
                    when others=>null;
                end case;
            end if;
        end if;
    end process;
    
    -- //****************************************************************************************************
    -- //  ģ������:50Mʱ�ӷ�Ƶ��1HZģ��
    -- //  ��������:
    -- //****************************************************************************************************
    process(clk,reset_n)
      begin 
        if(reset_n = '0')then
            clk_1hz <= '0';
            count <= "0000000000000000000000000";
        elsif(clk'event and clk = '1')then--�����ش���
            if(count = "1011111010111100001000000")then--
                count <= "0000000000000000000000000";
                clk_1hz <= not clk_1hz;
            else
                count <= count + '1';
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:�����ɨ��ʱ�Ӳ���ģ��
    -- //  ��������:
    -- //****************************************************************************************************
    process(clk,reset_n)
    begin
        if(reset_n = '0')then
            scan_count <= "00000000000000";
            clk_scan <= '0';
        elsif(clk'event and clk = '1')then--�����ش���
            if(scan_count = "10011100010000")then
                scan_count <= "00000000000000";
                clk_scan <= not clk_scan;
            else
                scan_count <= scan_count + '1';
            end if;
        end if;
    end process;
    process(clk_scan,reset_n)
    begin
        if(reset_n = '0')then
            seg_select <= "00";
        elsif(clk_scan'event and clk_scan = '1')then--�����ش���
            seg_select <= seg_select + '1';
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:�������ʾģ��
    -- //  ��������:
    -- //****************************************************************************************************
    process(reset_n,data_temp) 
    variable e,f,g:std_logic_vector(3 downto 0);  
    begin
        if(reset_n = '0')then
            data_temp_shi <= "0000";
            data_temp_ge <= "0000";
        else
            f := not data_temp(4 downto 1);
            g := "1010";
            e := "0000"; 
            for i in 15 downto 0 loop--���ü�������ʽ�����г�������
                if (f >= g) then 
                    f := f - g;
                    e := e + '1';
                else
                    exit; 
                end if; 
            end loop; 
            data_temp_shi <= e;
            data_temp_ge <= f;
        end if;
    end process; 
    
    process(clk)
    begin 
        if(clk'event and clk = '1')then--�����ش���
            case seg_select is
            when "00"=>--
                seg_wei <= "11111110";
                case (data_temp_ge) is
                    when "0000"=>seg_duan <= "11000000";--0
                    when "0001"=>seg_duan <= "11111001";--1
                    when "0010"=>seg_duan <= "10100100";--2
                    when "0011"=>seg_duan <= "10110000";--3
                    when "0100"=>seg_duan <= "10011001";--4
                    when "0101"=>seg_duan <= "10010010";--5
                    when "0110"=>seg_duan <= "10000010";--6
                    when "0111"=>seg_duan <= "11111000";--7
                    when "1000"=>seg_duan <= "10000000";--8
                    when "1001"=>seg_duan <= "10010000";--9
                    when others=>null;
                end case;
            when "01"=>--
                seg_wei <="11111101";
                case (data_temp_shi) is
                    when "0000"=>seg_duan <= "11000000";--0
                    when "0001"=>seg_duan <= "11111001";--1
                    when "0010"=>seg_duan <= "10100100";--2
                    when "0011"=>seg_duan <= "10110000";--3
                    when "0100"=>seg_duan <= "10011001";--4
                    when "0101"=>seg_duan <= "10010010";--5
                    when "0110"=>seg_duan <= "10000010";--6
                    when "0111"=>seg_duan <= "11111000";--7
                    when "1000"=>seg_duan <= "10000000";--8
                    when "1001"=>seg_duan <= "10010000";--9
                    when others=>null;
                end case;
            when others=>null;
            end case;
        end if;
    end process;
    
 end behave;
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
