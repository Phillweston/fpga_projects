/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� key.v
** �������ڣ�
** ������������������
** Ӳ��ƽ̨�������ϵ�һ�������� http://daxiguafpga.taobao.com
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module key(
           clk,
           key,
           key_out);
input clk;
input key; //ʱ�����룬��������
output key_out;//��������İ����ź����

wire clk;
wire key;

reg  key_out;

parameter s0=2'b00,s1=2'b01,s2=2'b10,s3=2'b11;
reg [1:0] state;

always @(posedge clk)
 begin
    case (state)
     s0:
      begin 
       key_out<=1'b1;
	   if(key==1'b0)
		  state<=s1;
	   else 
	      state<=s0;
	  end
	 s1:
	  begin 
	   if(key==1'b0)
		 state<=s2;
	   else 
	     state<=s0;
	   end 
	 s2:
	  begin 
	   if(key==1'b0)
		 state<=s3;
	   else 
	     state<=s0;    
	   end 
	 s3:
	   begin 
	    if(key==1'b0)
	     begin
		 key_out<=1'b0;
		 state<=s3;
		 end 
		else 
		 begin
		 key_out<=1'b1;
		 state<=s0;
	     end
	   end
	 default:
	     state<=s0;
    endcase
 end
endmodule

