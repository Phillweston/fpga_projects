----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:   
-- Design Name: 
-- Module Name:    plane - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--������ʾ����ʾ���ķɻ���״���ã�������ַ���0��ɵľ��Ƿɻ���ģ��
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity plane is
    port(
        y,x: in std_logic_vector(5 downto 0);----location of point��y����ĳһ�У�x����ĳһ�У����Ƕ�ά����
        data: out std_logic---yan se xin xi �ɻ�����ɫ�ź�
    );
end plane;

architecture Behavioral of plane is
    type rom_type is array(0 to 31) of std_logic_vector(31 downto 0);
    constant FONT: rom_type :=
    ("11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111111111111111111111",
     "11111111111111100111111111111111",
     "11111111111111100111111111111111",
     "11111111111111100111111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111110011001111111111111",
     "11111111111110011001111111111111",
     "11111111111110000001111111111111",
     "11111111111110000001111111111111",
     "11111111100000111100000111111111",
     "11111100000000100100000000111111",
     "11000000000000111100000000000011",
     "11000000000011000011000000000011",
     "11000001111111000011111110000011",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111111000011111111111111",
     "11111111111110000001111111111111",
     "11111111111100000000111111111111",
     "11111111110000100100001111111111",
     "11111111000000011000000011111111",
     "11111111111001111110011111111111",
     "11111111111111111111111111111111");

signal d:std_logic_vector(31 downto 0);
begin 

d<=FONT(conv_integer(y));
data<=not d(conv_integer(x));

end Behavioral;