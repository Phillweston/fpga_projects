//���ֲ���ģ��
module song(clk_6mhz,clk_4hz,speaker,high,med,low,k);    //ģ����Ϊsong���˿��б�
input clk_6mhz,clk_4hz; 
input k;                            //������������˿�
output speaker;                                      //����һ������˿�
output[3:0] high,med,low;                             
reg[3:0] high,med,low;                            //������3��4λ�Ĵ���
reg[13:0] divider,origin;                              //������2��14λ�Ĵ���
reg[9:0] counter;                                    //������1��10λ�Ĵ���
reg speaker;                                        
wire carry;
assign carry=(divider==16383);                         //������ֵ���
always @(posedge clk_6mhz)
    begin  if(carry) divider<=origin;
           else    divider<=divider+1;
    end
always @(posedge carry)
    begin speaker<=~speaker;
end                      //����Ƶ���������ź�
always @(posedge clk_4hz)
 begin
   case({high,med,low})                             //��Ƶ��Ԥ��
   'b000000000011:origin<=7281;                     //����3
   'b000000000101:origin<=8730;                     //����5
   'b000000000110:origin<=9565;                     //����6
   'b000000000111:origin<=10310;                    //����7
   'b000000010000:origin<=10647;                    //����1
   'b000000100000:origin<=11272;                    //����2
   'b000000110000:origin<=11831;                    //����3
   'b000001010000:origin<=12556;                    //����5
   'b000001100000:origin<=12974;                    //����6
   'b000001110000:origin<=13347;                    //����7
   'b000100000000:origin<=13516;                    //����1
   'b000000000000:origin<=16383;                    //��ֹ��
endcase
	
 end
always @(posedge clk_4hz)  
if (k==0) 
 begin
   if(counter==149)    counter<=0;                   //��ʱ����ʵ��ѭ������
   else               counter<=counter+1;
   case(counter)                                    //����
   0:  {high,med,low}<='b000000000011;              //����"3"
   1:  {high,med,low}<='b000000000011;              //����4��ʱ�ӽ���
   2:  {high,med,low}<='b000000000011;
   3:  {high,med,low}<='b000000000011;
   4:  {high,med,low}<='b000000000101;              //����"5"
   5:  {high,med,low}<='b000000000101;              //��3��ʱ�ӽ���
   6:  {high,med,low}<='b000000000101;
   7:  {high,med,low}<='b000000000110;              //����"6"
   8:  {high,med,low}<='b000000010000;              //����"1"
   9:  {high,med,low}<='b000000010000;              //��3��ʱ�ӽ���
   10: {high,med,low}<='b000000010000;
   11: {high,med,low}<='b000000100000;              //����"2"
   12: {high,med,low}<='b000000000110;              //����"6"
   13: {high,med,low}<='b000000010000;              //����"1"
   14: {high,med,low}<='b000000000101;              //����"5"
   15: {high,med,low}<='b000000000101;
   16: {high,med,low}<='b000001010000;              //����"5"
   17: {high,med,low}<='b000001010000;              //��3��ʱ�ӽ���
   18: {high,med,low}<='b000001010000;
   19: {high,med,low}<='b000100000000;              //����"1"
   20: {high,med,low}<='b000001100000;              //����"6"
   21: {high,med,low}<='b000001010000;              //����"5"
   22: {high,med,low}<='b000000110000;              //����"3"
   23: {high,med,low}<='b000001010000;              //����"5"
   24: {high,med,low}<='b000000100000;              //����"2"
   25: {high,med,low}<='b000000100000;              //����11��ʱ�ӽ���
   26: {high,med,low}<='b000000100000;
   27: {high,med,low}<='b000000100000;
   28: {high,med,low}<='b000000100000;
   29: {high,med,low}<='b000000100000;
   30: {high,med,low}<='b000000100000;
   31: {high,med,low}<='b000000100000;
   32: {high,med,low}<='b000000100000;
   33: {high,med,low}<='b000000100000;
   34: {high,med,low}<='b000000100000;
   35: {high,med,low}<='b000000110000;              //����"3"
   36: {high,med,low}<='b000000000111;              //����"7"
   37: {high,med,low}<='b000000000111;
   38: {high,med,low}<='b000000000110;              //����"6"
   39: {high,med,low}<='b000000000110;
   40: {high,med,low}<='b000000000101;              //����"5"
   41: {high,med,low}<='b000000000101;
   42: {high,med,low}<='b000000000101;
   43: {high,med,low}<='b000000000110;              //����"6"
   44: {high,med,low}<='b000000010000;              //����"1"
   45: {high,med,low}<='b000000010000;
   46: {high,med,low}<='b000000100000;              //����"2"
   47: {high,med,low}<='b000000100000;
   48: {high,med,low}<='b000000000011;              //����"3"
   49: {high,med,low}<='b000000000011;
   50: {high,med,low}<='b000000010000;              //����"1"
   51: {high,med,low}<='b000000010000;
   52: {high,med,low}<='b000000000110;              //����"6"
   53: {high,med,low}<='b000000000101;              //����"5"
   54: {high,med,low}<='b000000000110;              //����"6"
   55: {high,med,low}<='b000000010000;              //����"1"
   56: {high,med,low}<='b000000000101;              //����"5"
   57: {high,med,low}<='b000000000101;              //����8��ʱ�ӽ���
   58: {high,med,low}<='b000000000101;
   59: {high,med,low}<='b000000000101;
   60: {high,med,low}<='b000000000101;
   61: {high,med,low}<='b000000000101;
   62: {high,med,low}<='b000000000101;
   63: {high,med,low}<='b000000000101;
   64: {high,med,low}<='b000000110000;               //����"3"
   65: {high,med,low}<='b000000110000;               //��3��ʱ�ӽ���
   66: {high,med,low}<='b000000110000;
   67: {high,med,low}<='b000001010000;               //����"5"
   68: {high,med,low}<='b000000000111;               //����"7"
   69: {high,med,low}<='b000000000111;
   70: {high,med,low}<='b000000100000;               //����"2"
   71: {high,med,low}<='b000000100000;
   72: {high,med,low}<='b000000000110;               //����"6"
   73: {high,med,low}<='b000000010000;               //����"1"
   74: {high,med,low}<='b000000000101;               //����"5"
   75: {high,med,low}<='b000000000101;               //����4��ʱ�ӽ���
   76: {high,med,low}<='b000000000101;
   77: {high,med,low}<='b000000000101;
   78: {high,med,low}<='b000000000000;               //��ֹ��
   79: {high,med,low}<='b000000000000;
   80: {high,med,low}<='b000000000011;               //����"3"
   81: {high,med,low}<='b000000000101;               //����"5"
   82: {high,med,low}<='b000000000101; 
   83: {high,med,low}<='b000000000011;               //����"3"
   84: {high,med,low}<='b000000000101;               //����"5"
   85: {high,med,low}<='b000000000110;               //����"6"
   86: {high,med,low}<='b000000000111;               //����"7"
   87: {high,med,low}<='b000000100000;               //����"2"
   88: {high,med,low}<='b000000000110;               //����"6"
   89: {high,med,low}<='b000000000110;               //����6��ʱ�ӽ���
   90: {high,med,low}<='b000000000110;
   91: {high,med,low}<='b000000000110;
   92: {high,med,low}<='b000000000110;
   93: {high,med,low}<='b000000000110;
   94: {high,med,low}<='b000000000101;               //����"5"
   95: {high,med,low}<='b000000000110;               //����"6"
   96: {high,med,low}<='b000000010000;               //����"1"
   97: {high,med,low}<='b000000010000;               //��3��ʱ�ӽ���
   98: {high,med,low}<='b000000010000;
   99: {high,med,low}<='b000000100000;               //����"2"
   100: {high,med,low}<='b000001010000;              //����"5"
   101: {high,med,low}<='b000001010000;
   102: {high,med,low}<='b000000110000;              //����"3"
   103: {high,med,low}<='b000000110000;
   104: {high,med,low}<='b000000100000;              //����"2"
   105: {high,med,low}<='b000000100000;
   106: {high,med,low}<='b000000110000;              //����"3"
   107: {high,med,low}<='b000000100000;              //����"2"
   108: {high,med,low}<='b000000010000;              //����"1"
   109: {high,med,low}<='b000000010000;
   110: {high,med,low}<='b000000000110;              //����"6"
   111: {high,med,low}<='b000000000101;              //����"5"
   112: {high,med,low}<='b000000000011;              //����"3"
   113: {high,med,low}<='b000000000011;              //����4��ʱ�ӽ���
   114: {high,med,low}<='b000000000011;
   115: {high,med,low}<='b000000000011;
   116: {high,med,low}<='b000000010000;              //����"1"
   117: {high,med,low}<='b000000010000;              //����4��ʱ�ӽ���
   118: {high,med,low}<='b000000010000;
   119: {high,med,low}<='b000000010000;
   120: {high,med,low}<='b000000000110;              //����"6"
   121: {high,med,low}<='b000000010000;              //����"1"
   122: {high,med,low}<='b000000000110;              //����"6"
   123: {high,med,low}<='b000000000101;              //����"5"
   124: {high,med,low}<='b000000000011;              //����"3"
   125: {high,med,low}<='b000000000101;              //����"5"
   126: {high,med,low}<='b000000000110;              //����"6"
   127: {high,med,low}<='b000000010000;              //����"1"
   128: {high,med,low}<='b000000000101;              //����"5"
   129: {high,med,low}<='b000000000101;              //����6��ʱ�ӽ���
   130: {high,med,low}<='b000000000101;
   131: {high,med,low}<='b000000000101;
   132: {high,med,low}<='b000000000101;
   133: {high,med,low}<='b000000000101;
   134: {high,med,low}<='b000000110000;              //����"3"
   135: {high,med,low}<='b000001010000;              //����"5"
   136: {high,med,low}<='b000000100000;              //����"2"
   137: {high,med,low}<='b000000110000;              //����"3"
   138: {high,med,low}<='b000000100000;              //����"2"
   139: {high,med,low}<='b000000010000;              //����"1"
   140: {high,med,low}<='b000000000111;              //����"7"
   141: {high,med,low}<='b000000000111;
   142: {high,med,low}<='b000000000110;              //����"6"
   143: {high,med,low}<='b000000000110;
   144: {high,med,low}<='b000000000101;              //����"5"
   145: {high,med,low}<='b000000000101;              //����8��ʱ�ӽ���
   146: {high,med,low}<='b000000000101;
   147: {high,med,low}<='b000000000101;
   148: {high,med,low}<='b000000000101;
   149: {high,med,low}<='b000000000101;
   
   
endcase
end
else if( k==1)
begin
   if(counter==149)    counter<=0;                   //��ʱ����ʵ��ѭ������
   else               counter<=counter+1;
   case(counter)                                    //����
   0:  {high,med,low}<='b000000110000;              //����"3"
   1:  {high,med,low}<='b000000110000;              //����2��ʱ�ӽ���
   2:  {high,med,low}<='b000000100000;              //����2
   3:  {high,med,low}<='b000000100000;              //����2��ʱ�ӽ���
   4:  {high,med,low}<='b000000110000;              //����"3"
   5:  {high,med,low}<='b000000110000;              //��10��ʱ�ӽ���
   6:  {high,med,low}<='b000000110000;
   7:  {high,med,low}<='b000000110000;              
   8:  {high,med,low}<='b000000110000;             
   9:  {high,med,low}<='b000000110000;             
   10: {high,med,low}<='b000000110000;
   11: {high,med,low}<='b000000110000;             
   12: {high,med,low}<='b000000110000;              
   13: {high,med,low}<='b000000110000;         
   14: {high,med,low}<='b000000100000;              //����2
   15: {high,med,low}<='b000000100000;              //����2��ʱ�ӽ���
   16: {high,med,low}<='b000000110000;              //����"3"
   17: {high,med,low}<='b000000110000;              //��2��ʱ�ӽ���
   18: {high,med,low}<='b000000100000;              //����2
   19: {high,med,low}<='b000000100000;              //����2
   20: {high,med,low}<='b000000010000;              //����"1"
   21: {high,med,low}<='b000000010000;
   22: {high,med,low}<='b000000010000;
   23: {high,med,low}<='b000000010000;
   24: {high,med,low}<='b000000010000;
   25: {high,med,low}<='b000000010000;
   26: {high,med,low}<='b000000010000;
   27: {high,med,low}<='b000000010000;
   28: {high,med,low}<='b000000010000;
   29: {high,med,low}<='b000000010000;
   30: {high,med,low}<='b000000010000;
   31: {high,med,low}<='b000000010000;
   32: {high,med,low}<='b000000000110;//��6
   33: {high,med,low}<='b000000000110;
   34: {high,med,low}<='b000000010000;              //����"1"
   35: {high,med,low}<='b000000010000;              
   36: {high,med,low}<='b000000100000;              //��2  ��6��
   37: {high,med,low}<='b000000100000; 
   38: {high,med,low}<='b000000100000; 
   39: {high,med,low}<='b000000100000; 
   40: {high,med,low}<='b000000100000; 
   41: {high,med,low}<='b000000100000; 
   42: {high,med,low}<='b000000110000;               //����3
   43: {high,med,low}<='b000000110000;              
   44: {high,med,low}<='b000000100000;              //����"2"
   45: {high,med,low}<='b000000100000;
   46: {high,med,low}<='b000000010000;              //����"1"
   47: {high,med,low}<='b000000010000;
   48: {high,med,low}<='b000000000110;              //����"6"
   49: {high,med,low}<='b000000000110;
   50: {high,med,low}<='b000000010000;              //����"1"
   51: {high,med,low}<='b000000010000;
   52: {high,med,low}<='b000000000101;              //����"5"
   53: {high,med,low}<='b000000000101;              //����"5"
   54: {high,med,low}<='b000000000101; 
   55: {high,med,low}<='b000000000101; 
   56: {high,med,low}<='b000000000101;              //����"5"
   57: {high,med,low}<='b000000000101; 
   58: {high,med,low}<='b000000000101; 
   59: {high,med,low}<='b000000000101; 
   60: {high,med,low}<='b000000000101; 
   61: {high,med,low}<='b000000000101; 
   62: {high,med,low}<='b000000000101; 
   63: {high,med,low}<='b000000000101; 
   64: {high,med,low}<='b000000000101; 
   65: {high,med,low}<='b000000000101; 
66: {high,med,low}<='b000000000101; 
   67: {high,med,low}<='b000000000101; 
   68: {high,med,low}<='b000000110000;               //����"3"
   69: {high,med,low}<='b000000110000; 
   70: {high,med,low}<='b000000100000;               //����"2"
   71: {high,med,low}<='b000000100000;
   72: {high,med,low}<='b000000110000;               //����"3"
   73: {high,med,low}<='b000000110000;               //����"3"
   74: {high,med,low}<='b000000110000;               //����"3"
   75: {high,med,low}<='b000000110000;               //����"3"
   76: {high,med,low}<='b000000110000;               //����"3"
   77: {high,med,low}<='b000000110000;               //����"3"
   78: {high,med,low}<='b000000110000;               //����"3"
   79: {high,med,low}<='b000000110000;               //����"3"
   80: {high,med,low}<='b000000110000;               //����"3"
   81: {high,med,low}<='b000000110000;               //����"3"
   82: {high,med,low}<='b000000100000;               //����"2"
   83: {high,med,low}<='b000000100000;               
   84: {high,med,low}<='b000000110000;               //����"3"
   85: {high,med,low}<='b000000110000;               //����"3"
   86: {high,med,low}<='b000000100000;               //����"2"
   87: {high,med,low}<='b000000100000;               //����"2"
   88: {high,med,low}<='b000000010000;              //����"1"
   89: {high,med,low}<='b000000010000;              //����"1"
   90: {high,med,low}<='b000000010000;              //����"1"
   91: {high,med,low}<='b000000010000;              //����"1"
   92: {high,med,low}<='b000000010000;              //����"1"
   93: {high,med,low}<='b000000010000;              //����"1"
   94: {high,med,low}<='b000000010000;              //����"1"
   95: {high,med,low}<='b000000010000;              //����"1"
   96: {high,med,low}<='b000000010000;              //����"1"
   97: {high,med,low}<='b000000010000;              //����"1"
   98: {high,med,low}<='b000000010000;              //����"1"
   99: {high,med,low}<='b000000010000;              //����"1"
   100: {high,med,low}<='b000000010000;              //����"1"
   101: {high,med,low}<='b000000010000;              //����"1"
   102: {high,med,low}<='b000000010000;              //����"1"
   103: {high,med,low}<='b000000010000;              //����"1"
   104: {high,med,low}<='b000000010000;              //����"1"
   105: {high,med,low}<='b000000000110;              //����"6"
   106: {high,med,low}<='b000000000110;              //����"6"
   107: {high,med,low}<='b000000010000;              //����"1"
   108: {high,med,low}<='b000000010000;              //����"1"
   109: {high,med,low}<='b000000100000;               //����"2"
   110: {high,med,low}<='b000000100000;               //����"2"
   111: {high,med,low}<='b000000100000;               //����"2"
   112: {high,med,low}<='b000000100000;               //����"2"
   113: {high,med,low}<='b000000100000;               //����"2"
   114: {high,med,low}<='b000000100000;               //����"2"
   115: {high,med,low}<='b000000110000;               //����3
   116: {high,med,low}<='b000000110000;              
   117: {high,med,low}<='b000000100000;              //����"2"
   118: {high,med,low}<='b000000100000;
   119: {high,med,low}<='b000000010000;              //����"1"
   120: {high,med,low}<='b000000010000;
   121: {high,med,low}<='b000000000110;              //����"6"
   122: {high,med,low}<='b000000000110;
   123: {high,med,low}<='b000000010000;              //����"1"
   124: {high,med,low}<='b000000010000;
   125: {high,med,low}<='b000000100000;              //����"2"
   126: {high,med,low}<='b000000100000;              //����"2"
   127: {high,med,low}<='b000000100000;              //����"2"
   128: {high,med,low}<='b000000100000;              //����"2"
   129: {high,med,low}<='b000000100000;              //����"2"
   130: {high,med,low}<='b000000100000;              //����"2"
   131: {high,med,low}<='b000000100000;              //����"2"
   132: {high,med,low}<='b000000100000;              //����"2"
   133: {high,med,low}<='b000000100000;              //����"2"
   134: {high,med,low}<='b000000100000;              //����"2"
   135: {high,med,low}<='b000000100000;              //����"2"
   136: {high,med,low}<='b000000100000;              //����"2"
   137: {high,med,low}<='b000000100000;              //����"2"
   138: {high,med,low}<='b000000100000;              //����"2"
   139: {high,med,low}<='b000000100000;              //����"2"
   140: {high,med,low}<='b000000100000;              //����"2"
   141:  {high,med,low}<='b000000110000;              //����"3"
   142:  {high,med,low}<='b000000110000;              //����2��ʱ�ӽ���
   143:  {high,med,low}<='b000000100000;              //����2
   144:  {high,med,low}<='b000000100000;              //����2��ʱ�ӽ���
   145:  {high,med,low}<='b000000110000;              //����"3"
   146:  {high,med,low}<='b000000110000;              //��10��ʱ�ӽ���
   147:  {high,med,low}<='b000000110000;
   148:  {high,med,low}<='b000000110000;              
   149:  {high,med,low}<='b000000110000;  
  endcase
end
            
endmodule                                          //ģ��