/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� DDS.v
** �������ڣ�
** ����������DDS�źŷ�����Ƕ��ʽ�߼������ǵĵ���
** Ӳ��ƽ̨�������ϵ�һ�������� http://daxiguafpga.taobao.com
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module DDS(
           clk,
           reset_n,
           dds_data_out1,
           dds_data_out2,
           dds_data_out3
           );
input         clk;//ʱ������
input         reset_n;
output [9:0]  dds_data_out1;
output [9:0]  dds_data_out2;
output [9:0]  dds_data_out3;

wire          clk;
wire          reset_n;
wire    [9:0]  dds_data_out1;
wire    [9:0]  dds_data_out2;
wire    [9:0]  dds_data_out3;
//**************************************************//
//******************�����ز�1(500)**********************//
//**************************************************//
/**************������***************/
wire   [31:0] f32_bus1;//ACƵ�ʿ���������
wire   [9:0]  p_bus1;
wire   [31:0] reg32_out1;//32λ�Ĵ������
wire   [31:0] reg32_in1;//32λ�Ĵ�������
wire   [9:0]  reg10_in1;
wire   [9:0]  reg10_out_address1;
/************************************/

parameter [11:0] f32_bus_init1=12'd0;
parameter [9:0] p10_bus_init1=10'd0;//���ó�ʼ��λ

assign f32_bus1[31:20]=f32_bus_init1;//��ʼ��,��λ�õ�
assign f32_bus1[19:0]=20'd42950;//��λ��������DDS�����Ƶ��
assign p_bus1=p10_bus_init1;
/*********************Ԫ������************************************/
       adder_32 u1(.data1(f32_bus1),.data2(reg32_out1),.sum(reg32_in1));
       reg32    u2(.clk(clk),.reset_n(reset_n),.data_in(reg32_in1),.data_out(reg32_out1));
       adder_10 u3(.data1(p_bus1),.data2(reg32_out1[31:22]),.sum(reg10_in1));
       reg_10   u4(.clk(clk),.reset_n(reset_n),.data_in(reg10_in1),.data_out(reg10_out_address1));
       sin_rom  u5(.address(reg10_out_address1),.clock(clk),.q(dds_data_out1));//����
//**************************************************//
//******************�����ز�2(1K)**********************//
//**************************************************//
/**************������***************/
wire   [31:0] f32_bus2;//ACƵ�ʿ���������
wire   [9:0]  p_bus2;
wire   [31:0] reg32_out2;//32λ�Ĵ������
wire   [31:0] reg32_in2;//32λ�Ĵ�������
wire   [9:0]  reg10_in2;
wire   [9:0]  reg10_out_address2;
/************************************/

parameter [11:0] f32_bus_init2=12'd0;//
parameter [9:0] p10_bus_init2=10'd0;//���ó�ʼ��λ

assign f32_bus2[31:20]=f32_bus_init2;//��ʼ��,��λ�õ�
assign f32_bus2[19:0]=20'd85899;//��λ��������DDS�����Ƶ��
assign p_bus2=p10_bus_init2;
/*********************Ԫ������************************************/
       adder_32 u6(.data1(f32_bus2),.data2(reg32_out2),.sum(reg32_in2));
       reg32    u7(.clk(clk),.reset_n(reset_n),.data_in(reg32_in2),.data_out(reg32_out2));
       adder_10 u8(.data1(p_bus2),.data2(reg32_out2[31:22]),.sum(reg10_in2));
       reg_10   u9(.clk(clk),.reset_n(reset_n),.data_in(reg10_in2),.data_out(reg10_out_address2));
       sin_rom  u10(.address(reg10_out_address2),.clock(clk),.q(dds_data_out2));//����
//**************************************************//
//******************�����ز�3(1K,��λ��2�෴)**********************//
//**************************************************//
/**************������***************/
wire   [31:0] f32_bus3;//ACƵ�ʿ���������
wire   [9:0]  p_bus3;
wire   [31:0] reg32_out3;//32λ�Ĵ������
wire   [31:0] reg32_in3;//32λ�Ĵ�������
wire   [9:0]  reg10_in3;
wire   [9:0]  reg10_out_address3;
/************************************/

parameter [11:0] f32_bus_init3=12'd0;//
parameter [9:0] p10_bus_init3=10'd512;//���ó�ʼ��λ

assign f32_bus3[31:20]=f32_bus_init3;//��ʼ��,��λ�õ�
assign f32_bus3[19:0]=20'd85899;//��λ��������DDS�����Ƶ��
assign p_bus3=p10_bus_init3;
/*********************Ԫ������************************************/
       adder_32 u11(.data1(f32_bus3),.data2(reg32_out3),.sum(reg32_in3));
       reg32    u12(.clk(clk),.reset_n(reset_n),.data_in(reg32_in3),.data_out(reg32_out3));
       adder_10 u13(.data1(p_bus3),.data2(reg32_out3[31:22]),.sum(reg10_in3));
       reg_10   u14(.clk(clk),.reset_n(reset_n),.data_in(reg10_in3),.data_out(reg10_out_address3));
       sin_rom  u15(.address(reg10_out_address3),.clock(clk),.q(dds_data_out3));//����
endmodule





