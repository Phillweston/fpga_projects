// *******************************************************************************
// �����ļ�ģ��
// *******************************************************************************/
module fir_dac(
              clk,
              reset_n,
              key_in,
              sclk,                  //TLC5615 sclkʱ�ӽ�
              din,                   //TLC5615 din���ݽ�
              cs                    //TLC5615 csƬѡ
              );
input  clk;
input  reset_n;
input  key_in;
output sclk;
output din;
output cs;

wire [9:0]data_line;
wire [9:0]fir_data;
wire [9:0]data_in;
wire [9:0]fir_data_20;
fir fir_top(
           .clk(clk),
           .reset_n(reset_n),
           .data_in(data_in),  //г���ź�
           .fir_data(fir_data), //8�˲�֮����ź�
           .fir_data_20(fir_data_20)//21�˲�֮����ź�
           );
TLC5615 tlc5615_top(
           .clk(clk),//�ڲ�ʱ��
           .sclk(sclk),//TLC5615 sclkʱ�ӽ�
           .din(din),//TLC5615 din���ݽ�
           .cs(cs),//TLC5615 csƬѡ
           .din_in(data_line));//ʮλ�������� 
key key_top(
          .key_in(key_in),
          .data_out(data_line),
          .data1(fir_data),
          .data2(fir_data_20)
          );
endmodule
