/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� reg32.v
** �������ڣ�
** ��������:32λ�Ĵ���
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module reg32(
             clk,
             data_in,
             data_out);
input clk;
input [31:0] data_in;
output [31:0] data_out;

wire clk;
wire [31:0] data_in;
reg [31:0] data_out;

always @(posedge clk)
 begin
  data_out <= data_in;//�Ĵ�����
  end 
endmodule
