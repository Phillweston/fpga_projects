/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� reg_10.v
** ����������10λ�Ĵ���
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module reg_10(
             clk,
             data_in,
             data_out);
input clk;
input [8:0] data_in;
output [8:0] data_out;

wire clk;
wire [8:0] data_in;
reg [8:0] data_out;

always @(posedge clk)
 begin
  data_out<=data_in;//�Ĵ�����
  end 
endmodule