library IEEE;  
use IEEE.STD_LOGIC_1164.ALL;  
use IEEE.STD_LOGIC_ARITH.ALL;  
use IEEE.STD_LOGIC_UNSIGNED.ALL;  

entity ds18B20 is  
port(
    clk : in std_logic;---50MHz 
    rst_n: in std_logic; --��λ�ź�����
    one_wire  : inout std_logic;  --DS18B20������
    ---------------- 
    dataout : out std_logic_vector(7 downto 0); --������������
    en : out std_logic_vector(3 downto 0));  --�����λѡ�ź�  
end ds18B20;

architecture Behavioral of ds18B20 is  
signal dataout_buf:std_logic_vector(3 downto 0);   
signal count:std_logic_vector(17 downto 0); --��Ƶ������
signal cnt_scan:std_logic_vector(17 downto 0);   --����ܵ�ɨ����ʾ������
signal clk_1us:std_logic;-- 1MHz ʱ��

signal cnt_1us:integer range 0 to 750002;-- 1us��ʱ������
signal cnt_1us_clear:std_logic;-- ��1us��ʱ������
TYPE STATE_TYPE is (S00,S0,S1,S2,S3,S4,S5,S6,S7,
                    WRITE0,WRITE1,WRITE00,WRITE01,READ0,READ1,READ2,READ3);  --״̬��
signal state: STATE_TYPE;  --��ʼ״̬����Ϊ��λ״̬
signal one_wire_buf:std_logic;-- One-Wire���� ����Ĵ���
signal temperature_buf:std_logic_vector(15 downto 0);-- �ɼ������¶�ֵ��������δ����
signal DS18B20_DATA_buf:std_logic_vector(15 downto 0);-- �ɼ������¶�ֵ��������δ����
signal DS18B20_DATA_buf_temp:std_logic_vector(15 downto 0);-- �ɼ������¶�ֵ��������δ����
signal step:integer range 0 to 50;--��״̬�Ĵ��� 0~50
signal bit_valid:integer range 0 to 15;--��Чλ 
signal one_wire_in:std_logic;
signal t_buf:std_logic_vector(15 downto 0);
signal t_buf_temp:std_logic_vector(15 downto 0);
signal cnt:integer range 0 to 50;-- ������
-- //++++++++++++++++++++++++++++++++++++++
-- // ��Ƶ��50MHz->1MHz ��ʼ
-- //++++++++++++++++++++++++++++++++++++++
begin
    -- process (clk,rst_n)
    -- begin  
        -- if rising_edge(clk) then  
            -- if(rst_n='0') then  
                -- cnt <= 0;
            -- else
                -- if(cnt = 49)then
                  -- cnt <= 0;
                -- else
                  -- cnt <= cnt + 1;
                -- end if;
            -- end if;
        -- end if;
    -- end Process;  
      
    process (clk,rst_n)-- 1MHz ʱ��
    begin  
        if rising_edge(clk) then  
            if(rst_n='0') then  
                clk_1us <= '0';
            else
                if (cnt = 24)then
                  clk_1us <= not clk_1us;
                  cnt <= 0;
                else
                    cnt <= cnt + 1;
                  -- clk_1us <= '1';    
                end if;
            end if;
        end if;
    end Process;  
-- //--------------------------------------
-- // ��Ƶ��50MHz->1MHz ����
-- //--------------------------------------

-- //++++++++++++++++++++++++++++++++++++++
-- // ��ʱģ�� ��ʼ
-- //++++++++++++++++++++++++++++++++++++++
    process (clk_1us,cnt_1us_clear)-- 1MHz ʱ��
    begin  
        if rising_edge(clk_1us) then  
            if (cnt_1us_clear = '1')then
                cnt_1us <= 0;
            else
                cnt_1us <= cnt_1us + 1;
            end if;
        end if;
    end Process;
-- //--------------------------------------
-- // ��ʱģ�� ����
-- //--------------------------------------

-- //++++++++++++++++++++++++++++++++++++++
-- // DS18B20״̬�� ��ʼ
-- //++++++++++++++++++++++++++++++++++++++
-- //++++++++++++++++++++++++++++++++++++++
process (clk_1us,rst_n)-- 1MHz ʱ��
    begin  
        if rising_edge(clk_1us) then  
            if(rst_n='0') then  
                one_wire_buf <= 'Z';
                step         <= 0;
                state        <= S00;
            else
            case (state)is
            when S00=>              
                      temperature_buf <= "0000000000011111";
                      state           <= S0;
            when S0=>                    -- ��ʼ��
                      cnt_1us_clear <= '1';
                      one_wire_buf  <= '0';              
                      state         <= S1;
            when S1=>
                    cnt_1us_clear <= '0';
                    if (cnt_1us = 500)then         -- ��ʱ500us
                        cnt_1us_clear <= '1';
                        one_wire_buf  <= 'Z';  -- �ͷ�����
                        state         <= S2;
                    end if;
            when S2=>
                      cnt_1us_clear <= '0';
                      if (cnt_1us = 100)then         -- �ȴ�100us
                        cnt_1us_clear <= '1';
                        state         <= S3;
                      end if;
            when S3=>if (one_wire='0')then              -- ��18b20��������,��ʼ���ɹ�
                      state <= S4;
                    elsif (one_wire = '1')then          -- ����,��ʼ�����ɹ�,����S0
                      state <= S0;
                    end if;
            when S4=>
                      cnt_1us_clear <= '0';
                      if (cnt_1us = 400)then         -- ����ʱ400us
                        cnt_1us_clear <= '1';
                        state         <= S5;
                      end if;       
            when S5=>-- д����
                      if(step = 0)then       -- 0xCC
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 1)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 2)then             
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01; 
                      elsif (step = 3)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;                
                      elsif (step = 4)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 5)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 6)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 7)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 8)then-- 0x44
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 9)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 10)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 11)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 12)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 13)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 14)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 15)then
                        step  <= step + 1;
                        state <= WRITE0;
                      -- // ��һ��д��,750ms��,����S0
                      elsif (step = 16)then
                        one_wire_buf <= 'Z';
                        step         <= step + 1;
                        state        <= S6;                
                      -- // �ٴ�����0xCC��0xBE
                      elsif (step = 17)then-- 0xCC
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 18)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 19)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;                
                      elsif (step = 20)then
                        step  <= step + 1;
                        state <= WRITE01;
                        one_wire_buf <= '0';
                      elsif (step = 21)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 22)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 23)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 24)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;               
                      elsif (step = 25)then-- 0xBE
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 26)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;                
                      elsif (step = 27)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;                
                      elsif (step = 28)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;                
                      elsif (step = 29)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 30)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      elsif (step = 31)then
                        step  <= step + 1;
                        state <= WRITE0;
                      elsif (step = 32)then
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= WRITE01;
                      -- // �ڶ���д��,����S7,ֱ�ӿ�ʼ������
                      elsif (step = 33)then
                        step  <= step + 1;
                        state <= S7;
                      end if;
            when S6=>
                      cnt_1us_clear <= '0';
                      if (cnt_1us = 750000 or one_wire='1')then     -- ��ʱ750ms!!!!
                        cnt_1us_clear <= '1';
                        state         <= S0;    -- ����S0,�ٴγ�ʼ��
                      end if;
            when S7=>                     -- ������
                      if(step = 34)then
                        bit_valid    <= 0;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;
                      elsif (step = 35)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;
                      elsif (step = 36)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;
                      elsif (step = 37)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;               
                      elsif (step = 38)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 39)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;               
                      elsif (step = 40)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 41)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;
                      elsif (step = 42)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 43)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;
                      elsif (step = 44)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      else if (step = 45)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 46)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 47)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 48)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 49)then
                        bit_valid    <= bit_valid + 1;
                        one_wire_buf <= '0';
                        step         <= step + 1;
                        state        <= READ0;                
                      elsif (step = 50)then
                        step  <= 0;
                        state <= S0;
                      end if;
                     end if;
				when WRITE0=>
                      cnt_1us_clear <= '0';
                      one_wire_buf  <= '0';-- ���0             
                      if (cnt_1us = 80)then-- ��ʱ80us
                        cnt_1us_clear <= '1';
                        one_wire_buf  <= 'Z'; -- �ͷ����ߣ��Զ�����                
                        state<= WRITE00;
                      end if;
				when WRITE00=>
						state <= S5;
				when WRITE01=>-- ��״̬
						state <= WRITE1;
				when WRITE1=>
						cnt_1us_clear <= '0';
                      one_wire_buf  <= 'Z';    -- ���1   �ͷ����ߣ��Զ�����
                      if (cnt_1us = 80)then        -- ��ʱ80us
                        cnt_1us_clear <= '1';
                        state<= S5; 
                       end if;
				when READ0=>state <= READ1;-- ����ʱ״̬
				when READ1=>
                      cnt_1us_clear <= '0';
                      one_wire_buf  <= 'Z';    -- �ͷ�����
                      if (cnt_1us = 10)then       -- ����ʱ10us
                        cnt_1us_clear <= '1';
                        state<= READ2;
                    end if;
				when READ2=>-- ��ȡ����
                      temperature_buf(bit_valid) <= one_wire;
                      state<= READ3;
				when READ3=>
                      cnt_1us_clear <= '0';
                      if (cnt_1us = 55)then-- ����ʱ55us
                        cnt_1us_clear <= '1';
                        state<= S7;
                    end if;
				when others=> state<=S00;
            end case;
		end if;
     end if;
end process;

    one_wire <= one_wire_buf;         -- ע��˫��ڵ�ʹ��
-- //--------------------------------------
-- // DS18B20״̬�� ����
-- //--------------------------------------
-- //++++++++++++++++++++++++++++++++++++++
-- // �Բɼ������¶Ƚ��д��� ��ʼ
-- //++++++++++++++++++++++++++++++++++++++
    process (temperature_buf)
    begin  
        t_buf <= temperature_buf and "0000011111111111";--07FF;
    end Process;  
-- //--------------------------------------
-- // �Բɼ������¶Ƚ��д������
-- //--------------------------------------
process (clk,rst_n)
begin
    if rising_edge(clk) then  
        if(rst_n='0')then
            DS18B20_DATA_buf <="0000000000000000";
            DS18B20_DATA_buf_temp <="0000000000000000";
            -- //��λ��ȫ������
        else
          t_buf_temp <= t_buf;
          DS18B20_DATA_buf_temp(15 downto 0) <=CONV_STD_LOGIC_VECTOR((CONV_INTEGER(t_buf(3 downto 0)) * 10),16);-- С�����һλ
          DS18B20_DATA_buf(3 downto 0) <= DS18B20_DATA_buf_temp(7 downto 4);
          
          if(t_buf_temp(7 downto 4) >= "1010")then -- ��λ
            DS18B20_DATA_buf(7 downto 4)   <= t_buf(7 downto 4) - "1010";
          else
            DS18B20_DATA_buf(7 downto 4)   <= t_buf(7 downto 4);   
          end if;
          
          if(t_buf_temp(7 downto 4) >= "1010")then -- ʮλ
            DS18B20_DATA_buf(11 downto 8)   <= t_buf(11 downto 8) + "0001";
          else
            DS18B20_DATA_buf(11 downto 8)   <= t_buf(11 downto 8);
          end if;
       -- // DS18B20_DATA_buf[15:12] = temperature_buf[12] ? 1 : 0;  
       -- // ��������ʾ�������Ǹ����ġ��������������� 
        end if;
    end if;
end Process;
-- //////////////////////////////////////////////////////////////////////////////////////////////////
-- //��Ƶ������
process (clk,rst_n)
begin
    if rising_edge(clk) then  
        if(rst_n='0')then
        count<="000000000000000000";	
        else
            count<=count+'1';
      -- //���������������Ŀ����Ϊ������ʾ����ܵ�  ʮλ  ��λ  С����  С�����һλ  ͬ��
      -- //������������������ʾɨ��Ҳ�õ���һ��λ��ļ�������
        end if;
    end if;
end Process;

process (clk)
begin
    if rising_edge(clk) then 
      case (count(17 downto 16))is
      -- //  Ҳ�Ƿ�Ƶ�Ĺؼ�
      -- //  ͨ����������Ƶ������ͬʱ�����ڣ���ʾ�¶ȵ�ʮλ  ��λ  С����  С�����һλ
      when "00"=> dataout_buf<=DS18B20_DATA_buf(3 downto 0);  --//С�����һλ  
      when "01"=> dataout_buf<="1010";                --//С���� 
      when "10"=> dataout_buf<=DS18B20_DATA_buf(7 downto 4);  --//��λ 
      when "11"=> dataout_buf<=DS18B20_DATA_buf(11 downto 8); --//ʮλ 
      end case;
    end if;
end Process;
-- //��Ƶ������
process (clk,rst_n)
begin
    if rising_edge(clk)then  
        if(rst_n='0')then
            cnt_scan<="000000000000000000";
        else
            cnt_scan<=cnt_scan+'1';
-- //���������������Ŀ����Ϊ������ʾ����ܵ�  ʮλ  ��λ  С����  С�����һλ�Ͷ�ȡDS18B20���¶�ֵͬ��
-- //�����������ʱ�εĶ�ȡDS18B20���¶�ֵҲ�õ���һ��λ��ļ�������
        end if;
    end if;
end Process;

process(cnt_scan)
begin
   case(cnt_scan(17 downto 16))is
                -- //case���Ĺ����ǰ����������������
                -- //�޸�cnt_scan[17:16]�������޸�����ܵ���ʾƵ�ʡ�
       when "00"=>
          en <= "1110";  --//������һλ����� .��ʾС�������һλ
       when "01"=>
          en <= "1101";  --//�����ڶ�λ����� ����������Ŀ������ʾ С����
       when "10"=>
          en <= "1101";  --//�����ڶ�λ����� ����������Ŀ������ʾ ��λ
       when "11"=>
          en <= "1011";  --//��������λ����� ������ʾ ʮλ
       when others=>
          en <= "1111";  --//�����ڰ�λ�����
    end case;
end Process;

process(dataout_buf)
begin
	case(dataout_buf)is
		when "0000"=>
			dataout<="11000000"; --//�����������ʾ0�Ķ���
		when "0001"=>
			dataout<="11111001"; --//�����������ʾ1�Ķ���
		when "0010"=>
			dataout<="10100100"; --//�����������ʾ2�Ķ���
		when "0011"=>
			dataout<="10110000"; --//�����������ʾ3�Ķ���
		when "0100"=>
			dataout<="10011001"; --//�����������ʾ4�Ķ���
		when "0101"=>
			dataout<="10010010"; --//�����������ʾ5�Ķ���
		when "0110"=>
			dataout<="10000010"; --//�����������ʾ6�Ķ���
		when "0111"=>
			dataout<="11111000"; --//�����������ʾ7�Ķ���
		when "1000"=>
			dataout<="11000000"; --//�����������ʾ8�Ķ���
		when "1001"=>
			dataout<="10010000"; --//�����������ʾ9�Ķ���	
		when "1010"=>
			dataout<="01111111"; --//�����������ʾС����Ķ���
		when others=>
			dataout<="10000000";
	 end case;
end Process;
end Behavioral; 



