/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ�TLC615.v
** �������ڣ�2012.10.10
** ����������ʹ��10λ����DAоƬTLC5615�������ź�ת��Ϊģ���źţ�������DAоƬVDD=5V,VREF=3.3V 
             ���㹫ʽ��Vout=VREF*(N/1024) NΪ10λ��������
** �������̣����������ڳ���ı�10λ������������DAоƬ��Vout�������Ӧ��ѹ
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module TLC5615
       (clk,                   //�ڲ�ʱ��
        sclk,                  //TLC5615 sclkʱ�ӽ�
        din,                   //TLC5615 din���ݽ�
        cs,                    //TLC5615 csƬѡ
        din_in);               //ʮλ�������� 
            
input      clk;
input [9:0]din_in;
output     din;
output     cs;
output     sclk;

reg        din;
reg        cs;
reg        sclk;
reg [3:0]  count1,count2,count3;
reg [9:0]  din_reg;                //10λ���ݼĴ���
initial                          //��ʼ��
begin
  cs=1;
  din=0;
  count1=0;
  count2=0;
  count3=0;
//  din_reg=10'b00_0000_1111;                    //ʵ���߿��Ը�����Ҫ�޸�10Ϊ��������
end

/************************************************/
/*** sclk��Ƶ������Ϊ5MHz ***/
always@(posedge clk)
begin
  if(count3==4'd9)
  begin   
     sclk<=~sclk;
     count3<=0;
  end
  else
    count3<=count3+1'b1;
end
/*********��DDS���������ݽ��мĴ�**********/
always@(posedge clk)
  begin
   din_reg<=din_in;
  end

 
/*** TLC5615 csƬѡ ***/
always@(negedge sclk)
begin
  if(count1>=4'd12&&count1<4'd15)
  begin
     cs<=1;                                      //����Ƭѡ
     count1<=count1+4'd1;
  end
  else if(count1==4'd15)
  begin
    count1<=0;
  end
  else
  begin
    cs<=0;                                       //����Ƭѡ
    count1<=count1+4'd1;
  end 
end 

/*** 10λ�������������ģת��������12λ���ͷ�ʽ��10λ��Чλ+2λ���λ�� ***/
always@(posedge sclk)
begin
  if(cs==0)
  begin
  case(count2)
  4'd0:din<=1'd0;                                //��Чλ
  
  4'd1:begin din<=din_reg[9];end                 //10λ��Чλ      
  4'd2:begin din<=din_reg[8];end
  4'd3:begin din<=din_reg[7];end 
  4'd4:begin din<=din_reg[6];end 
  4'd5:begin din<=din_reg[5];end 
  4'd6:begin din<=din_reg[4];end 
  4'd7:begin din<=din_reg[3];end 
  4'd8:begin din<=din_reg[2];end 
  4'd9:begin din<=din_reg[1];end
  4'd10:begin din<=din_reg[0];end 
  
  4'd11:begin din<=1'd0;end                      //���λ ��0����
  4'd12:begin din<=1'd0;end                      //���λ ��0����
  
  4'd13:din<=1'd0;                               //��Чλ
  4'd14:din<=1'd0;                               //��Чλ
  4'd15:din<=1'd0;                               //��Чλ
  default:begin count2<=0;din<=0;end
  endcase
  end
  if(count2==4'd15)
   count2<=0;
  else
   count2<=count2+4'd1;
end 

endmodule 
  