-- ******************************************************************************
-- ����ģ��
-- ��������
-- �ϵ����Ȱ���key5�������и�λ����
-- (1)����key3���������һ�����룬�������һ���������key3������ڶ������룬�ڶ�������������ɺ����key3��
--      ������������룬����������������ɺ����key3��������ĸ����룬���ĸ�����������ɺ����key3��������ɣ�
-- (2)ֻ������������ȷ����ܽ����޸����룻
-- (3)�޸�����������£�
        -- ����key1�����޸�����״̬��Ȼ��ͨ��key2����ѡ�񰴼���ÿ����һ�����룬����key3����һ�Σ������������һλ��������һ�����룬
        -- 4������������ɺ���key4������ȷ�����������ͻ�����װ�ؽ�ȥ������λ����ܻ���ʾ��ǰ���������Ĵ���
        -- ȡ���޸����밴��key5��
-- *******************************************************************************
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
entity control is
port(
    clk:in std_logic;                               --50Mʱ������
    reset_n:in std_logic;                           --��λ�ź�����
    set_signal:in std_logic;                        --�������밴��
    select_signal:in std_logic;                     --
    ok_signal:in std_logic;                         --
    set_ok_signal:in std_logic;                         --
    
    fm_time_over:in std_logic;                      --������20����Ӧ����ź�
    fm_20:in std_logic;
    password1_out:out std_logic_vector(3 downto 0); --
    password2_out:out std_logic_vector(3 downto 0); --
    password3_out:out std_logic_vector(3 downto 0); --
    password4_out:out std_logic_vector(3 downto 0); --
    ok_signal_counter_out:out std_logic_vector(2 downto 0);--�ĸ�����ܵı��
    motor_open:out std_logic;                       --������ر�־
    start_flag:out std_logic;
    password_yes:out std_logic;
    password_no:out std_logic;
    password_set_out:out std_logic
);
end control;
architecture control_behave of control is 
signal key_counter:std_logic_vector(3 downto 0);    --�������´���������
signal password_set:std_logic;                      --���������־����1��Ϊ�������룬��0��Ϊû����������
signal password_set_finish:std_logic;               --�������óɹ��ź�
signal ok_signal_counter:std_logic_vector(2 downto 0);--�����������������
signal current_password1:std_logic_vector(3 downto 0);--��ǰ��һ������
signal current_password2:std_logic_vector(3 downto 0);--��ǰ�ڶ�������
signal current_password3:std_logic_vector(3 downto 0);--��ǰ����������
signal current_password4:std_logic_vector(3 downto 0);--��ǰ���ĸ�����
signal current_password1_temp:std_logic_vector(3 downto 0);--��ǰ��һ������
signal current_password2_temp:std_logic_vector(3 downto 0);--��ǰ�ڶ�������
signal current_password3_temp:std_logic_vector(3 downto 0);--��ǰ����������
signal current_password4_temp:std_logic_vector(3 downto 0);--��ǰ���ĸ�����
signal password1:std_logic_vector(3 downto 0);      --�����һ������
signal password2:std_logic_vector(3 downto 0);      --����ڶ�������
signal password3:std_logic_vector(3 downto 0);      --�������������
signal password4:std_logic_vector(3 downto 0);      --������ĸ�����
signal set_signal_re1:std_logic;
signal set_signal_re2:std_logic;
signal password_yes_temp:std_logic;
signal password_no_temp:std_logic;
signal start_flag_reg:std_logic;
type state is(
            prepare,--׼��״̬
            start--��ʼ״̬
            );
signal current_state:state;--һ��ʼ����׼��״̬

type set_state is(
            prepare,--׼��״̬
            start--��ʼ״̬
            );
signal current_set_state:set_state;--һ��ʼ����׼��״̬
begin
    password_set_out <= not password_set;
    ok_signal_counter_out <= ok_signal_counter;
    start_flag <= start_flag_reg;
    -- //****************************************************************************************************
    -- //  ģ������:�������������ź�password_set
    -- //  ��������:
    -- //****************************************************************************************************
    process(clk,reset_n)
    begin
        if(reset_n = '0')then
            password_set <= '0';
            current_set_state <= prepare;
            
            current_password1 <= "0001";
            current_password2 <= "0001";
            current_password3 <= "0001";
            current_password4 <= "0001";
            
        elsif(clk'event and clk = '0')then--�½��ش���
            if((password_yes_temp = '1'and password_no_temp = '0') or password_set = '1')then--ֻ������������ȷ������޸�����
                case current_set_state is
                when prepare=>
                    if(set_signal = '0')then
                        current_set_state <= start;
                        password_set <= '1';
                    else
                        current_set_state <= prepare;
                        password_set <= '0';
                    end if;
                when start =>
                    if(set_ok_signal = '0')then--�������
                        --����װ������
                        current_password1 <= current_password1_temp;
                        current_password2 <= current_password2_temp;
                        current_password3 <= current_password3_temp;
                        current_password4 <= current_password4_temp;
                        current_set_state <= prepare;
                        password_set <= '0';
                    else
                        password_set <= '1';
                        current_set_state <= start;
                    end if;
                when others=>null;
                end case;
            else
                null;
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:Υʱ�źŵĲ���
    -- //  ��������:
    -- //****************************************************************************************************
    process(clk,reset_n)
    begin
        if(reset_n = '0')then
            current_state <= prepare; 
            start_flag_reg <= '0';
        elsif(clk'event and clk = '1')then--�������ش���
            if(password_set = '0')then--����������״̬
                case current_state is
                when prepare=>
                    if(select_signal = '0')then
                        start_flag_reg <= '1';
                        current_state <= start; 
                    else
                        start_flag_reg <= '0';
                        current_state <= prepare;
                    end if;
                when start=>
                    if(ok_signal_counter = "100")then--�����������
                        start_flag_reg <= '0';
                        current_state <= prepare;
                    elsif(fm_time_over = '1')then--��������Ӧ20s���
                        start_flag_reg <= '0';
                        current_state <= prepare; 
                    else--����δ���
                        start_flag_reg <= '1';
                        current_state <= start; 
                    end if;
                end case;
            else
                current_state <= prepare; 
                start_flag_reg <= '0';
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:����������������
    -- //  ��������:
    -- //****************************************************************************************************
    process(select_signal,reset_n)
    begin
        if(reset_n = '0')then
            key_counter <= "0000";
        elsif(select_signal'event and select_signal = '0')then--�½��ش���
            if(key_counter = "1001")then
                key_counter <= "0000";
            else
                key_counter <= key_counter + '1';
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:ͳ����������ĸ���4��
    -- //  ��������:
    -- //****************************************************************************************************
    process(ok_signal,reset_n)
    begin
        if(reset_n = '0')then
            ok_signal_counter <= "000";
        elsif(ok_signal'event and ok_signal = '0')then--�½��ش���
            if(fm_20 = '0')then--�ڲ�Υʱ������¿��Խ�����������
                if(ok_signal_counter = "100")then
                    ok_signal_counter <= "001";
                    --�����������
                else
                    ok_signal_counter <= ok_signal_counter + '1';
                end if;
            else
                ok_signal_counter <= "000";
            end if;
        end if;
    end process;
    -- //****************************************************************************************************
    -- //  ģ������:�洢��������ĸ���4��
    -- //  ��������:
    -- //****************************************************************************************************
    process(clk,reset_n)
    begin
        if(reset_n = '0')then
        ----------------------------------
            current_password1_temp <= "0000";
            current_password2_temp <= "0000";
            current_password3_temp <= "0000";
            current_password4_temp <= "0000";
        ----------------------------------
            password_yes_temp <= '0';
            password_no_temp <= '1';
            password1 <= "0000";
            password2 <= "0000";
            password3 <= "0000";
            password4 <= "0000";
            motor_open <= '1';--�����
        elsif(clk'event and clk = '1')then--�����ش���
            if(fm_20 = '0')then--�ڲ�Υʱ������¿��Խ�����������
                case ok_signal_counter is
                when "001"=>
                            if(password_set = '0')then--����������
                                password1 <= key_counter;
                            else--��������
                                current_password1_temp <= key_counter;
                                password1 <= "0000";
                                motor_open <= '1';--�����
                                password_yes_temp <= '0';
                                password_no_temp <= '0';
                            end if;
                when "010"=>
                            if(password_set = '0')then--����������
                                password2 <= key_counter;
                            else--��������
                                current_password2_temp <= key_counter;
                                password2 <= "0000";
                                motor_open <= '1';--�����
                                password_yes_temp <= '0';
                                password_no_temp <= '0';
                            end if;
                when "011"=>
                            if(password_set = '0')then--����������
                                password3 <= key_counter;
                            else--��������
                                current_password3_temp <= key_counter;
                                password3 <= "0000";
                                motor_open <= '1';--�����
                                password_yes_temp <= '0';
                                password_no_temp <= '0';
                            end if;
                when "100"=>
                            if(password_set = '0')then--����������
                                password4 <= key_counter;
                                if(current_password1 = password1 and 
                                    current_password2 = password2 and 
                                        current_password3 = password3 and 
                                            current_password4 = password4)then
                                    password_yes_temp <= '1';
                                    password_no_temp <= '0';
                                    motor_open <= '0';--�����
                                else
                                    password_yes_temp <= '0';
                                    password_no_temp <= '1';
                                    motor_open <= '1';--�����
                                end if;
                            else--��������
                                current_password4_temp <= key_counter;
                                password4 <= "0000";
                                motor_open <= '1';--�����
                                password_yes_temp <= '0';
                                password_no_temp <= '0';
                            end if;
                when others=>null;
                end case;
            else
                password_yes_temp <= '0';
                password_no_temp <= '1';
                password1 <= "0000";
                password2 <= "0000";
                password3 <= "0000";
                password4 <= "0000";
                motor_open <= '1';--�����
            end if;
        end if;
    end process;
    -- ��������������״̬ʱ���������ǲ�����
    password_yes <= not ((password_yes_temp) and (not password_set));--����ɫled��141����
    password_no <= not ((password_no_temp) and (not password_set));--�Ӻ�ɫled��142����
    
    -- //****************************************************************************************************
    -- //  ģ������:�������ʾ����ѡ��ģ��
    -- //  ��������:
    -- //****************************************************************************************************
    process(reset_n,password_set,
    current_password1_temp,current_password2_temp,current_password3_temp,current_password4_temp,
    password1,password2,password3,password4)
    begin
        if(reset_n = '0')then
            password1_out <= "0000";
            password2_out <= "0000";
            password3_out <= "0000";
            password4_out <= "0000";
        elsif(password_set = '1')then--��������
            password1_out <= current_password1_temp;
            password2_out <= current_password2_temp;
            password3_out <= current_password3_temp;
            password4_out <= current_password4_temp;
        else--����������
            password1_out <= password1;
            password2_out <= password2;
            password3_out <= password3;
            password4_out <= password4;
        end if;
    end process;
    

end control_behave;












