-- ��1��miso �C ���豸�������룬���豸���������
-- ��2��mosi �C ���豸������������豸�������룻
-- ��3��SCLK �C ʱ���źţ������豸������
-- ��4��CS �C ���豸ʹ���źţ������豸���ơ�
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity spi_out is
port(
     clk_in:in std_logic;   --ʱ������ 50M
     miso:in std_logic;     --���ź�
     cs:out std_logic;      --Ƭѡ�ź�
     mosi:out std_logic;    --���ź�
     sck_out:out std_logic;  --ʱ���ź�
     received_data_out:out std_logic_vector(7 downto 0)
);
end spi_out;
architecture spi_behave of spi_out is
signal data_out:std_logic_vector(7 downto 0);--���͵�8bit����
signal num:     integer range 0 to 9;       --������
signal clk_div: std_logic;                  --��Ƶ
signal gain_data:std_logic_vector(8 downto 0);
begin 
   sck_out<=clk_div;
   data_out<="01100110";--Ԥ�跢������
   -- *************************************************
   -- ʱ�ӷ�Ƶģ�飬��50Mʱ�ӽ��з�Ƶ��Ȼ�󽫷�Ƶ���ʱ����Ϊ
   -- spi��ʱ���źţ���Ƶ���ʱ���ź�Ϊ5M
   -- *************************************************
   process(clk_in)--��Ƶ
    variable counter:integer range 0 to 4;
     begin 
        if(clk_in'event and clk_in='1')then
           if(counter=4)then 
                counter:=0;
                clk_div<=not clk_div;
           else 
                counter:=counter+1;
           end if;
        end if;
   end process;
   -- *************************************************
   -- ���ݷ���ģ��
   -- ��num��1~8�ķ�Χ�ڽ�8bit�����ݽ��з��ͣ����͵�ͬʱ
   -- cs�ڵ͵�ƽ��ʱ����Ч��ѡͨspi�Ĵӻ�
   -- *************************************************
   process(clk_div)--����,�½���
      begin
        if(clk_div'event and clk_div='0')then 
            if(num=9)then-- ��numΪ9��ʱ���num�������㣬�Խ�����һ�����ݷ���
                num<=0;
            else 
                num<=num+1;
            end if;
            if(num>0 and num<9)then--��num��1~8�ķ�Χ�ڽ�8bit�����ݽ��з���
               cs<='0';--cs�ڵ͵�ƽ��ʱ����Ч��ѡͨspi�Ĵӻ�
               mosi<=data_out(8-num);--��num�������½�8bit����������ͳ�ȥ����λ��ǰ����λ�ں�
            else 
               cs<='1';--������ɺ󣬽�cs���ߣ���ѡͨspi�ӻ�
               mosi<='Z';--���͸���̬�ź�
            end if;
        end if;
   end process;
   

   process(clk_div)
      variable num:integer range 0 to 9;
      begin 
          if(clk_div'event and clk_div='1')then 
                if(num>0 and num<9)then 
				  gain_data(9-num)<=miso;
                  num:=num+1;
                  if(num = 8)then
                    received_data_out<=gain_data(7 downto 0);
                  end if;
                elsif(num=9)then
                  num:=0;
                else
				  num:=num+1;
                end if;
		  end if;
		  
   end process;
end  spi_behave; 
   
   
   
   
   
   
   
         
         
         
   
   
   
   
   
                