/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� reg32.v
** �������ڣ�
** ��������:32λ�Ĵ���
** Ӳ��ƽ̨�������ϵ�һ��������
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module reg32(clk,reset_n,data_in,data_out);
input clk;
input reset_n;
input [31:0] data_in;
output [31:0] data_out;

wire clk;
wire reset_n;
wire [31:0] data_in;
reg [31:0] data_out;

always @(posedge clk or negedge reset_n)
 begin
  if(!reset_n)
   data_out<=32'd0;
  else
   data_out<=data_in;
  end 
endmodule
